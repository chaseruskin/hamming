--------------------------------------------------------------------------------
--! Project  : crus.ecc.hamming
--! Engineer : Chase Ruskin
--! Created  : 2022-10-02
--! Entity   : hamming_ecc
--! Details  :
--!     @todo: write general overview of component and its behavior
--!
--------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

entity hamming_ecc is 

    -- @todo: define port interface

end entity hamming_ecc;


architecture rtl of hamming_ecc is

    -- @todo: define internal signals/components

begin

    -- @todo: describe the circuit

end architecture rtl;
