-- Testbench for the `hamm_dec` module using file IO and event logging.

library ieee;
use ieee.std_logic_1164.all;

library test;
use test.verb.all;

library std;
use std.textio.all;

library work;
use work.hamm_pkg.all;

entity hamm_dec_tb is 
    generic (
        --! number of parity bits to decode (excluding 0th DED bit)
        PARITY_BITS : positive range 2 to positive'high := 4 
    );
end entity hamm_dec_tb;


architecture sim of hamm_dec_tb is

    -- This record is automatically @generated by Verb.
    -- It is not intended for manual editing.
    type hamm_dec_bfm is record
        encoding: logics(block_size(PARITY_BITS)-1 downto 0);
        message: logics(data_size(PARITY_BITS)-1 downto 0);
        corrected: logic;
        valid: logic;
    end record;

    signal bfm: hamm_dec_bfm;

    --! internal testbench signals
    constant DELAY : time := 10 ns;
    signal halt: boolean := false;

    file events: text open write_mode is "events.log";

begin

    dut: entity work.hamm_dec
    generic map (
        PARITY_BITS => PARITY_BITS
    ) port map (
        encoding  => bfm.encoding,
        message   => bfm.message,
        corrected => bfm.corrected,
        valid     => bfm.valid
    );

    --! assert the received outputs match expected model values
    bench: process
        file inputs  : text open read_mode is "inputs.txt";
        file outputs : text open read_mode is "outputs.txt";

        -- This procedure is automatically @generated by Verb.
        -- It is not intended for manual editing.
        procedure send(file i: text) is
            variable row: line;
        begin
            if endfile(i) = false then
                readline(i, row);
                drive(row, bfm.encoding);
            end if;
        end procedure;

        -- This procedure is automatically @generated by Verb.
        -- It is not intended for manual editing.
        procedure compare(file e: text; file o: text) is
            variable row: line;
            variable mdl: hamm_dec_bfm;
        begin
            if endfile(o) = false then
                readline(o, row);
                load(row, mdl.message);
                assert_eq(e, bfm.message, mdl.message, "message");
                load(row, mdl.corrected);
                assert_eq(e, bfm.corrected, mdl.corrected, "corrected");
                load(row, mdl.valid);
                assert_eq(e, bfm.valid, mdl.valid, "valid");
            end if;
        end procedure;
    begin
        -- @todo: drive UUT and check circuit behavior
        while not endfile(inputs) loop
            --! read given inputs from file
            send(inputs);

            wait for DELAY;

            compare(events, outputs);
        end loop;
        complete(events, halt);
    end process;

end architecture;