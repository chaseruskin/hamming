-- Testbench for the `hamm_enc` module using file IO and event logging.

library ieee;
use ieee.std_logic_1164.all;

library work;
use work.hamm_pkg.all;

library test;
use test.verb.all;

library std;
use std.textio.all;

entity hamm_enc_tb is 
    generic (
        PARITY_BITS : positive range 2 to positive'high := 4
    );
end entity hamm_enc_tb;


architecture sim of hamm_enc_tb is

    -- This record is automatically @generated by Verb.
    -- It is not intended for manual editing.
    type hamm_enc_bfm is record
        message: logics(data_size(PARITY_BITS)-1 downto 0);
        encoding: logics(block_size(PARITY_BITS)-1 downto 0);
    end record;
    
    signal bfm: hamm_enc_bfm;

    --! internal testbench signals
    constant DELAY: time := 10 ns;
    signal halt: boolean := false;

    file events: text open write_mode is "events.log";
begin

    dut: entity work.hamm_enc
        generic map (
            PARITY_BITS => PARITY_BITS
        ) port map (
            message   => bfm.message,
            encoding  => bfm.encoding
        );

    --! assert the received outputs match expected model values
    bench: process
        file inputs  : text open read_mode is "inputs.txt";
        file outputs : text open read_mode is "outputs.txt";

        -- This procedure is automatically @generated by Verb.
        -- It is not intended for manual editing.
        procedure send(file i: text) is
            variable row: line;
        begin
            if endfile(i) = false then
                readline(i, row);
                drive(row, bfm.message);
            end if;
        end procedure;

        -- This procedure is automatically @generated by Verb.
        -- It is not intended for manual editing.
        procedure compare(file e: text; file o: text) is
            variable row: line;
            variable mdl: hamm_enc_bfm;
        begin
            if endfile(o) = false then
                readline(o, row);
                load(row, mdl.encoding);
                assert_eq(e, bfm.encoding, mdl.encoding, "encoding");
            end if;
        end procedure;
    begin
        while not endfile(inputs) loop
            send(inputs);
            wait for DELAY;
            compare(events, outputs);
        end loop;
        complete(events, halt);
    end process;

end architecture sim;